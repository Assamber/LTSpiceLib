*Mar 22, 2010
*Doc. ID: 90302, Rev. A
*File Name: part irf9640_sihf9640_PS.txt and part irf9640_sihf9640_PS.spi
*This document is intended as a SPICE modeling guideline and does not
*constitute a commercial product datasheet. Designers should refer to the
*appropriate data sheet of the same number for guaranteed specification
*limits.
.SUBCKT irf9640 1 2 3
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*Commercial Use or Resale Restricted *
*   by Symmetry License Agreement    *
**************************************
* Model generated on May 21, 96
* Model format: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
* Default values used in MM:
* The voltage-dependent capacitances are
* not included. Other default values are:
*   RS=0 RD=0 LD=0 CBD=0 CBS=0 CGBO=0
.MODEL MM PMOS LEVEL=1 IS=1e-32
+VTO=-3.8062 LAMBDA=0.0228396 KP=10.7224
+CGSO=1.09465e-05 CGDO=1e-11
RS 8 3 0.101556
D1 1 3 MD
.MODEL MD D IS=1e-17 RS=0.185714 N=1.5 BV=200
+IBV=0.00025 EG=1.2 XTI=4 TT=1e-07
+CJO=1.22255e-09 VJ=2.42988 M=0.605683 FC=0.493595
RDS 3 1 2e+06
RD 9 1 0.261579
RG 2 7 6.81119
D2 5 4 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=8.6947e-10 VJ=2.34088 M=0.9 FC=1e-08
D3 5 0 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=1e-10 N=0.402798 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 1.8148e-09
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 6 0 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=1e-10 N=0.402798
.ENDS

