* DIODES INCORPORATED AND ITS AFFILIATED COMPANIES AND SUBSIDIARIES (COLLECTIVELY, "DIODES") 
* PROVIDE THESE SPICE MODELS AND DATA (COLLECTIVELY, THE "SM DATA") "AS IS" AND WITHOUT ANY 
* REPRESENTATIONS OR WARRANTIES, EXPRESS OR IMPLIED, INCLUDING ANY WARRANTY OF MERCHANTABILITY 
* OR FITNESS FOR A PARTICULAR PURPOSE, ANY WARRANTY ARISING FROM COURSE OF DEALING OR COURSE OF 
* PERFORMANCE, OR ANY WARRANTY THAT ACCESS TO OR OPERATION OF THE SM DATA WILL BE UNINTERRUPTED, 
* OR THAT THE SM DATA OR ANY SIMULATION USING THE SM DATA WILL BE ERROR FREE. TO THE MAXIMUM 
* EXTENT PERMITTED BY LAW, IN NO EVENT WILL DIODES BE LIABLE FOR ANY DIRECT OR INDIRECT, 
* SPECIAL, INCIDENTAL, PUNITIVE OR CONSEQUENTIAL DAMAGES ARISING OUT OF OR IN CONNECTION WITH 
* THE PRODUCTION OR USE OF SM DATA, HOWEVER CAUSED AND UNDER WHATEVER CAUSE OF ACTION OR THEORY 
* OF LIABILITY BROUGHT (INCLUDING, WITHOUT LIMITATION, UNDER ANY CONTRACT, NEGLIGENCE OR OTHER 
* TORT THEORY OF LIABILITY), EVEN IF DIODES HAS BEEN ADVISED OF THE POSSIBILITY OF SUCH DAMAGES, 
* AND DIODES' TOTAL LIABILITY (WHETHER IN CONTRACT, TORT OR OTHERWISE) WITH REGARD TO THE SM 
* DATA WILL NOT, IN THE AGGREGATE, EXCEED ANY SUMS PAID BY YOU TO DIODES FOR THE SM DATA.



*ZETEX ZVN0545A Spice Model v1.0 Last Revised 20/5/04
    *
    *
    .SUBCKT ZVN0545A 3 4 5
    *                D G S
    M1 6 20 8 8 MOSMOD
    M2 6 20 8 8 MOSMODS
    RG 4 2 55
    RIN 2 8 200E6
    RD 3 6 RMOD1 40
    RS 8 5 RMOD1 2.5 
    RL 3 5 200E6
    C1 2 8 160E-12
    C2 17 3 2E-12 
    D1 5 3 DMOD1
    D2 17 3 DMOD2
    Egs1 2 17 2 8 1
    Egt1 2 20 21 5 1
    Vgt1 5 22 1
    Igt1 5 21 1
    Rgt 21 22 RMOD2 1
    .MODEL MOSMOD NMOS VTO=2.26 IS=1E-15 KP=.59 CBD=15E-12 PB=1 LAMBDA=4.9E-3
    .MODEL MOSMODS NMOS VTO=1.9 IS=1E-15 KP=0.02 PB=1
    .MODEL DMOD1 D IS=2E-13 RS=10 N=1.01 IKF=3e-3
    .MODEL DMOD2 D CJO=25e-12 IS=1e-30 N=10
    .MODEL RMOD1 RES (TC1=8E-3 TC2=1.7E-5)
    .MODEL RMOD2 RES (TC1=-2.5e-3 TC2=3.3e-6)
    .ENDS
    *
    *$
    *