***************************************************************												
*	Infineon	Technologies	AG									
*	GUMMEL-POON	MODEL	IN	SPICE	2G6	SYNTAX				
*	VALID	UP	TO	10	GHZ							
*	>>>	BFR360F	<<<								
*	(C)	2019	Infineon	Technologies	AG							
*	Version	1.0	January 2019							
***************************************************************			
.OPTION GMIN= 1.00e-12
*BFR360F C B E
.SUBCKT BFR360F 1 2 3

CBEPAR 22 33 5.287E-14
CBCPAR 22 11 3.004E-13
CCEPAR 11 33 1.51929E-13
LB   22 20 2.93767E-10
LE   33 30 3.6E-10
RCI 11 10 0.0009993
CBEPCK 20 30  5.29743E-15
CCEPCK 10 30  5.7E-14
CBCPCK 20 10  1.589E-15
LBX    20 2 1.2E-10
LEX    30 3 1.2E-10
LCX    10 1 2E-10


Q1 11 22 33 M_BFR360F

.MODEL 	M_BFR360F	NPN(	
+	TNOM	=	25									
+	IS	=	9.721E-17									
+	BF	=	170.4									
+	NF	=	0.999									
+	VAF	=	49.37									
+	IKF	=	0.3647									
+	ISE	=	4.419E-15									
+	NE	=	1.999									
+	BR	=	10.36		
+	NR	=	0.9996		
+	VAR	=	2.773	
+	IKR	=	0.03687		
+	ISC	=	3.261E-16		
+	NC	=	1.34		
+	RB	=	6		
+	IRB	=	1E-05		
+	RBM	=	2	
+	RE	=	0.4105		
+	RC	=	8.385	
+	XTB	=	-0.1945		
+	EG	=	1.11		
+	XTI	=	5.65		
+	CJE	=	4.2E-13		
+	VJE	=	0.631654		
+	MJE	=	0.247368		
+	TF	=	8.7E-12		
+	XTF	=	97.8956		
+	VTF	=	0.742		
+	ITF	=	0.695		
+	PTF	=	5		
+	CJC	=	7.071E-14		
+	VJC	=	0.774619		
+	MJC	=	0.846923		
+	XCJC	=	0.7499		
+	TR	=	7.927E-09
+	CJS	=	6.05859E-15		
+	MJS	=	2.12235
+   VJS =   0.272069 		
+	FC	=	0.63		
+	KF	=	2E-10		
+	AF	=	2)
***************************************************************					
					

.ENDS BFR360F
