* DIODES INCORPORATED AND ITS AFFILIATED COMPANIES AND SUBSIDIARIES (COLLECTIVELY, "DIODES") 
* PROVIDE THESE SPICE MODELS AND DATA (COLLECTIVELY, THE "SM DATA") "AS IS" AND WITHOUT ANY 
* REPRESENTATIONS OR WARRANTIES, EXPRESS OR IMPLIED, INCLUDING ANY WARRANTY OF MERCHANTABILITY 
* OR FITNESS FOR A PARTICULAR PURPOSE, ANY WARRANTY ARISING FROM COURSE OF DEALING OR COURSE OF 
* PERFORMANCE, OR ANY WARRANTY THAT ACCESS TO OR OPERATION OF THE SM DATA WILL BE UNINTERRUPTED, 
* OR THAT THE SM DATA OR ANY SIMULATION USING THE SM DATA WILL BE ERROR FREE. TO THE MAXIMUM 
* EXTENT PERMITTED BY LAW, IN NO EVENT WILL DIODES BE LIABLE FOR ANY DIRECT OR INDIRECT, 
* SPECIAL, INCIDENTAL, PUNITIVE OR CONSEQUENTIAL DAMAGES ARISING OUT OF OR IN CONNECTION WITH 
* THE PRODUCTION OR USE OF SM DATA, HOWEVER CAUSED AND UNDER WHATEVER CAUSE OF ACTION OR THEORY 
* OF LIABILITY BROUGHT (INCLUDING, WITHOUT LIMITATION, UNDER ANY CONTRACT, NEGLIGENCE OR OTHER 
* TORT THEORY OF LIABILITY), EVEN IF DIODES HAS BEEN ADVISED OF THE POSSIBILITY OF SUCH DAMAGES, 
* AND DIODES' TOTAL LIABILITY (WHETHER IN CONTRACT, TORT OR OTHERWISE) WITH REGARD TO THE SM 
* DATA WILL NOT, IN THE AGGREGATE, EXCEED ANY SUMS PAID BY YOU TO DIODES FOR THE SM DATA.

*---------- DMP510DL Spice Model ----------
.SUBCKT DMP510DL 10 20 30 
*     TERMINALS:  D  G  S
M1 1 2 3 3 PMOS L = 1E-006 W = 1E-006 
RD 10 1 1.961 
RS 30 3 0.001 
RG 20 2 916 
CGS 2 3 2.2E-011 
EGD 12 30 2 1 1 
VFB 14 30 0 
FFB 2 1 VFB 1 
CGD 13 14 3.8E-011 
R1 13 30 1 
D1 13 12 DLIM 
DDG 14 15 DCGD 
R2 12 15 1 
D2 30 15 DLIM 
DSD 10 3 DSUB 
.MODEL PMOS PMOS LEVEL = 3 U0 = 400 VMAX = 1E+006 ETA = 0.001 
+ TOX = 6E-008 NSUB = 1E+016 KP = 0.2606 KAPPA = 49.86 VTO = -1.522 
.MODEL DCGD D CJO = 6.69E-012 VJ = 1 M = 0.1 
.MODEL DSUB D IS = 9.14E-010 N = 1.637 RS = 0.1748 BV = 66.94 CJO = 1E-015 VJ = 0.1 M = 0.1851 
.MODEL DLIM D IS = 0.0001 
.ENDS
*Diodes DMP510DL Spice Model v1.0 Last Revised 2015/9/24